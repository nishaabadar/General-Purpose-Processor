LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY decod IS
	PORT (s  : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			En : IN STD_LOGIC ;
			y 	: OUT STD_LOGIC_VECTOR(15 downto 0)) ;
END decod;

ARCHITECTURE Behaviour OF decod IS
	SIGNAL Ens : STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN
Ens <= En & s(3) & s(2)&s(1)&s(0);
WITH Ens SELECT
	y <=  "1000000000000000" WHEN "10000",--0
			"0100000000000000" WHEN "10001",--1
			"0010000000000000" WHEN "10010",--2
			"0001000000000000" WHEN "10011",--3
			"0000100000000000" WHEN "10100",--4
			"0000010000000000" WHEN "10101",--5
			"0000001000000000" WHEN "10110",--6
			"0000000100000000" WHEN "10111",--7
			"0000000010000000" WHEN "11000",--8
			"0000000000000000" WHEN OTHERS;
END Behaviour;

	